library ieee;
use ieee.std_logic_1164.all;
use std.numeric_std.all;





entity I2C_controllerNew is



end entity;






architecture rtl of I2C_controllerNew is




begin






end architecture;